module 4b5b_encoder;


endmodule
